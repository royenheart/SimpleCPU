`define PipInitStage 2'b00   //流水线初始阶段
`define PipInStage 2'b01     //流水线写入阶段
`define PipKeepStage 2'b10   //流水线保持阶段
`define PipOutStage 2'b11    //流水线写出阶段
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/03/06 19:37:32
// Design Name: 
// Module Name: ALU_test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ALU_test(

    );

    reg [4:0] opt;
    reg [31:0] in_1;
    reg [31:0] in_2;
    wire [31:0] out;
    wire zero;
    ALU alu1(.op(opt),.A(in_1),.B(in_2),.out(out),.zero(zero));
    initial begin
            opt = 5'b00000;
            in_1 = 108;
            in_2 = 62;
        #20 in_1 = 32'h80000074;
            in_2 = 32'h80000079;
        #20 in_1 = 32'h80000074;
            in_2 = 200;
        #20 in_1 = 32'h80000074;
            in_2 = 62;
            
       #20     opt = 5'b00001;
            in_1 = 32'hf2340000;
            in_2 = 32'h80000000;
        #20 in_1 = 32'h7fffffff;
            in_2 = 32'h70000001;
        #20 in_1 = 32'hffffffff;
            in_2 = 32'h00000001;
        #20 in_1 = 32'hf1a2c371;
            in_2 = 32'h7230ff45;


        #20 opt = 5'b000010;
            in_1 = 32'h0000006c;
            in_2 = 32'h0000003e;
        #20 in_1 = 32'h0000003e;
            in_2 = 32'h0000006c;
        #20 in_1 = 32'h0000006c;
            in_2 = 32'h8000003e;
        #20 in_1 = 32'h8000006c;
            in_2 = 32'h8000003e;
            
       #20     opt = 5'b00011;
            in_1 = 32'hf2340000;
            in_2 = 32'h80000000;
        #20 in_1 = 32'h7fffffff;
            in_2 = 32'h70000001;
        #20 in_1 = 32'hffffffff;
            in_2 = 32'h00000001;
        #20 in_1 = 32'hf1a2c371;
            in_2 = 32'h7230ff45;
            
        //AND
        #20 opt = 5'b00100;
            in_1 = 32'h72340000;
            in_2 = 32'h60000000;
        #20 in_1 = 32'h7fffffff;
            in_2 = 32'h00000000;

        //OR
        #20 opt = 5'b00101;
            in_1 = 32'h00000000;
            in_2 = 32'h00000000;
        #20 in_1 = 32'h7fffffff;
            in_2 = 32'hf0000001;
        
        //XOR
        #20 opt = 5'b00110;
            in_1 = 32'ha0000000;
            in_2 = 32'h50000000;
        #20 in_1 = 32'h7fffffff;
            in_2 = 32'hf0000001;

        #20 opt = 5'b00111;
            in_1 = 32'ha0000000;
            in_2 = 32'h50000000;
        #20 in_1 = 32'h7fffffff;
            in_2 = 32'hf0000001;
                
                
        #20 opt = 5'b01000;
            in_1 = 32'ha0000000;
            in_2 = 32'h50000000;
        #20 in_1 = 32'h7fffffff;
            in_2 = 32'hf0000001;
        #20 in_1 = 108;
            in_2 = 62;
        #20 in_1 = 62;
            in_2 = 32'h07234000;
        #20 in_1 = 32'hf0000001;
            in_2 = -62;
        #20 in_1 = -62;
            in_2 = -108;
               
               
        #20 opt = 5'b01001;
            in_1 = 32'ha0000000;
            in_2 = 32'h50000000;
        #20 in_1 = 32'h7fffffff;
            in_2 = 32'hf0000001;
               
                   
        //SAL
        #20 opt = 5'b01010;
            in_1 = 32'h7234abcc;
            in_2 = 32'h00000010;
        #20 in_1 = 32'h7230ff45;
            in_2 = 32'h00000016;
        #20 in_1 = 32'hf0001231;
            in_2 = 32'h00000020;
        #20 in_1 = 32'hf1a2c371;
            in_2 = 32'h00000009;
            
        //SAR
        #20 opt = 5'b01011;
            in_1 = 32'h7234abcc;
            in_2 = 32'h00000010;
        #20 in_1 = 32'h7230ff45;
            in_2 = 32'h00000016;
        #20 in_1 = 32'hf0001231;
            in_2 = 32'h00000020;
        #20 in_1 = 32'hf1a2c371;
            in_2 = 32'h00000009;
            
        #20 opt = 5'b01100;
            in_1 = 32'h7234abcc;
            in_2 = 32'h00000010;
        #20 in_1 = 32'h7230ff45;
            in_2 = 32'h00000016;
        #20 in_1 = 32'hf0001231;
            in_2 = 32'h00000020;
        #20 in_1 = 32'hf1a2c371;
            in_2 = 32'h00000009;


        #20 opt = 5'b01101;
            in_1 = 32'h7234abcc;
            in_2 = 32'h7234abcc;
        #20 in_1 = 32'h7230ff45;
            in_2 = 32'h00000016;
        #20 in_1 = 32'hf0001231;
            in_2 = 32'hf0001231;
            
        #20 opt = 5'b01110;
            in_1 = 32'h7234abcc;
            in_2 = 32'h7234abcc;
        #20 in_1 = 32'h7230ff45;
            in_2 = 32'h00000016;
        #20 in_1 = 32'hf0001231;
            in_2 = 32'hf0001231;
            
    end 
endmodule